`timescale 1 ns / 1 ps

module Read_weightnbais_TB ();

//************************Do Not Remove************************//
	initial begin
		$dumpfile("Read_weightnbais_TB.vcd");
		$dumpvars();
	end
//*************************************************************//

reg [15:0]t0,t1,t2,t3,t4;
reg [15:0]c1_w[0:5][0:0][4:0][4:0];
reg [15:0]c1_b[0:5];
reg [15:0]c3_w[0:15][5:0][4:0][4:0];
reg [15:0]c3_b[0:15];

initial begin
	#0
	$readmemh ("D:/FYP/FYP/weights/c1_weight.txt", c1_w);
    $readmemh ("D:/FYP/FYP/weights/c1_bias.txt", c1_b);
    $readmemh ("D:/FYP/FYP/weights/c3_weight.txt", c3_w);
    $readmemh ("D:/FYP/FYP/weights/c3_bias.txt", c3_b);
	t0 = 0;
	t1 = 0;
	t2 = 0;
	t3 = 0;
	t4 = 0;
	//c1_w*************
	#1
	t0 = c1_w[0][0][0][0];
	t1 = c1_w[0][0][1][1];
	t2 = c1_w[0][0][2][2];
	t3 = c1_w[0][0][3][3];
	t4 = c1_w[0][0][4][4];
	#1
	t0 = c1_w[1][0][0][0];
	t1 = c1_w[1][0][1][1];
	t2 = c1_w[1][0][2][2];
	t3 = c1_w[1][0][3][3];
	t4 = c1_w[1][0][4][4];
	#1
	t0 = c1_w[5][0][0][0];
	t1 = c1_w[5][0][1][1];
	t2 = c1_w[5][0][2][2];
	t3 = c1_w[5][0][3][3];
	t4 = c1_w[5][0][4][4];
	//***********************

	//c1_b*****************
	#1
	t0 = c1_b[0];
	t1 = c1_b[1];
	t2 = c1_b[3];
	t3 = c1_b[4];
	t4 = c1_b[5];
	//************************

	//c3_w*****************
	#1
	t0 = c3_w[0][0][0][0];
	t1 = c3_w[0][0][1][1];
	t2 = c3_w[0][0][2][2];
	t3 = c3_w[0][0][3][3];
	t4 = c3_w[0][0][4][4];
	#1
	t0 = c3_w[0][5][0][0];
	t1 = c3_w[0][5][1][1];
	t2 = c3_w[0][5][2][2];
	t3 = c3_w[0][5][3][3];
	t4 = c3_w[0][5][4][4];
	#1
	t0 = c3_w[1][0][0][0];
	t1 = c3_w[1][0][1][1];
	t2 = c3_w[1][0][2][2];
	t3 = c3_w[1][0][3][3];
	t4 = c3_w[1][0][4][4];	
	#1
	t0 = c3_w[1][5][0][0];
	t1 = c3_w[1][5][1][1];
	t2 = c3_w[1][5][2][2];
	t3 = c3_w[1][5][3][3];
	t4 = c3_w[1][5][4][4];
	#1
	t0 = c3_w[15][0][0][0];
	t1 = c3_w[15][0][1][1];
	t2 = c3_w[15][0][2][2];
	t3 = c3_w[15][0][3][3];
	t4 = c3_w[15][0][4][4];	
	#1
	t0 = c3_w[15][5][0][0];
	t1 = c3_w[15][5][1][1];
	t2 = c3_w[15][5][2][2];
	t3 = c3_w[15][5][3][3];
	t4 = c3_w[15][5][4][4];
	//************************

	//c3_b*****************
	#1
	t0 = c3_b[0];
	t1 = c3_b[4];
	t2 = c3_b[8];
	t3 = c3_b[11];
	t4 = c3_b[15];
	//************************

	#1
	$finish();
end

endmodule

