`timescale 1 ns / 1 ps

module Read_WB (


);



endmodule  
